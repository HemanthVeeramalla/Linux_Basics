#or gate
module or_gate(out,a,b);
input a,b;
output out;
assign out=a|b;
endmodule
